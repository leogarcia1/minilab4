`include "systolic_array_tc.svh"

module memA_tb();

