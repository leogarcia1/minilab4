`include "systolic_array_tc.svh"

module memB_tb();

